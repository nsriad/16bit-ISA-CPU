//=============================================
// Global Definitions for 16-bit ISA CPU
//=============================================
`define WORD_WIDTH 16
`define REG_COUNT  8
